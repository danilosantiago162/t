CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1610 30 100 10
176 80 1364 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 1 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
62
13 Logic Switch~
5 266 2043 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -17 7 -9
3 V18
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3277 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 252 1912 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -17 7 -9
3 V17
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4212 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 184 1794 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4720 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 183 1741 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V15
-9 -30 12 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5551 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 182 1684 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -17 7 -9
3 V14
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6986 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 165 1451 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8745 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 162 1327 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9592 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 868 1078 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8748 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 860 958 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7168 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 150 1119 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
631 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 143 1046 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9466 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 139 980 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3266 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 136 913 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7693 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 142 784 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3723 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 142 676 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3440 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 139 586 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6263 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 142 281 0 1 11
0 41
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4900 0 0
2
5.9012e-315 0
0
13 Logic Switch~
5 137 144 0 1 11
0 43
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8783 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 628 1980 0 3 22
0 6 7 5
0
0 0 624 0
4 7400
-7 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
3221 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 506 1921 0 3 22
0 2 3 6
0
0 0 624 0
4 7400
-7 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
3215 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 732 1933 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7903 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 371 1973 0 3 22
0 2 4 3
0
0 0 624 0
4 7400
-7 -24 21 -16
4 U11D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
7121 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 517 2034 0 3 22
0 3 4 7
0
0 0 624 0
4 7400
-7 -24 21 -16
4 U11C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
4484 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 441 1698 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
5.9012e-315 0
0
5 7409~
219 354 1723 0 3 22
0 12 10 8
0
0 0 624 0
6 74LS09
-21 -24 21 -16
4 U12A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
7804 0 0
2
5.9012e-315 0
0
8 2-In OR~
219 247 1762 0 3 22
0 9 11 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5523 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 608 1329 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 525 1356 0 3 22
0 14 15 13
0
0 0 624 0
4 7400
-7 -24 21 -16
4 U11B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3465 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 452 1426 0 3 22
0 16 17 15
0
0 0 624 0
4 7400
-7 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
8396 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 330 1464 0 3 22
0 18 18 17
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U8D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
3685 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 326 1314 0 3 22
0 19 18 14
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
7849 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 328 1388 0 3 22
0 19 19 16
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
6343 0 0
2
5.9012e-315 0
0
6 74266~
219 970 1020 0 3 22
0 23 22 20
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
7376 0 0
2
5.9012e-315 0
0
6 74266~
219 397 989 0 3 22
0 28 27 21
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
9156 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 1058 998 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 614 962 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
5.9012e-315 0
0
8 3-In OR~
219 533 989 0 4 22
0 26 21 25 24
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
4459 0 0
2
5.9012e-315 0
0
9 2-In AND~
219 275 1037 0 3 22
0 31 30 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3760 0 0
2
5.9012e-315 0
0
9 2-In AND~
219 273 904 0 3 22
0 32 29 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
754 0 0
2
5.9012e-315 0
0
5 7405~
219 220 1028 0 2 22
0 30 31
0
0 0 624 0
6 74LS05
-21 -24 21 -16
3 U9B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 6 0
65 0 0 0 6 2 9 0
1 U
9767 0 0
2
5.9012e-315 0
0
5 7405~
219 219 895 0 2 22
0 29 32
0
0 0 624 0
6 74LS05
-21 -24 21 -16
3 U9A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 6 0
65 0 0 0 6 1 9 0
1 U
7978 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 743 695 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3142 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 666 721 0 3 22
0 36 35 33
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3284 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 289 775 0 3 22
0 37 34 35
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
659 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 450 680 0 3 22
0 38 39 36
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3800 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 288 595 0 3 22
0 37 37 38
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6792 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 621 460 0 1 2
10 40
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 618 395 0 1 2
10 42
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6316 0 0
2
5.9012e-315 0
0
9 Inverter~
13 497 479 0 2 22
0 41 40
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 7 0
1 U
8734 0 0
2
5.9012e-315 0
0
9 Inverter~
13 495 415 0 2 22
0 43 42
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
7988 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 614 338 0 1 2
10 44
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3217 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 606 268 0 1 2
10 45
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3965 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 600 207 0 1 2
10 46
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8239 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 598 148 0 1 2
10 47
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
828 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 593 94 0 1 2
10 48
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6187 0 0
2
5.9012e-315 0
0
14 Logic Display~
6 592 19 0 1 2
10 49
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7107 0 0
2
5.9012e-315 0
0
6 74266~
219 486 347 0 3 22
0 43 41 44
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
6433 0 0
2
5.9012e-315 0
0
9 2-In XOR~
219 492 277 0 3 22
0 43 41 45
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
8559 0 0
2
5.9012e-315 0
0
5 7433~
219 486 214 0 3 22
0 43 41 46
0
0 0 624 0
6 74LS33
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 2 3 1 2 3 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3674 0 0
2
5.9012e-315 0
0
8 2-In OR~
219 486 162 0 3 22
0 43 41 47
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5697 0 0
2
5.9012e-315 0
0
10 2-In NAND~
219 494 106 0 3 22
0 43 41 48
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3805 0 0
2
5.9012e-315 0
0
9 2-In AND~
219 493 45 0 3 22
0 43 41 49
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5219 0 0
2
5.9012e-315 0
0
73
1 1 2 0 0 4224 0 2 20 0 0 2
264 1912
482 1912
3 2 3 0 0 4096 0 22 20 0 0 4
398 1973
458 1973
458 1930
482 1930
0 2 4 0 0 12432 0 0 23 8 0 2
339 2043
493 2043
3 1 3 0 0 4224 0 22 23 0 0 4
398 1973
465 1973
465 2025
493 2025
3 1 5 0 0 4224 0 19 21 0 0 3
655 1980
732 1980
732 1951
3 1 6 0 0 4224 0 20 19 0 0 4
533 1921
582 1921
582 1971
604 1971
3 2 7 0 0 4224 0 23 19 0 0 4
544 2034
582 2034
582 1989
604 1989
1 2 4 0 0 128 0 1 22 0 0 4
278 2043
339 2043
339 1982
347 1982
1 1 2 0 0 128 0 2 22 0 0 4
264 1912
339 1912
339 1964
347 1964
3 1 8 0 0 4224 0 25 24 0 0 3
375 1723
441 1723
441 1716
1 1 9 0 0 4224 0 4 26 0 0 4
195 1741
226 1741
226 1753
234 1753
3 2 10 0 0 4224 0 26 25 0 0 4
280 1762
317 1762
317 1732
330 1732
1 2 11 0 0 4224 0 3 26 0 0 4
196 1794
226 1794
226 1771
234 1771
1 1 12 0 0 4224 0 5 25 0 0 4
194 1684
322 1684
322 1714
330 1714
3 1 13 0 0 4224 0 28 27 0 0 3
552 1356
608 1356
608 1347
3 1 14 0 0 4224 0 31 28 0 0 4
353 1314
493 1314
493 1347
501 1347
3 2 15 0 0 8320 0 29 28 0 0 4
479 1426
493 1426
493 1365
501 1365
3 1 16 0 0 4224 0 32 29 0 0 4
355 1388
420 1388
420 1417
428 1417
3 2 17 0 0 4224 0 30 29 0 0 4
357 1464
420 1464
420 1435
428 1435
1 2 18 0 0 12288 0 6 30 0 0 4
177 1451
181 1451
181 1473
306 1473
1 1 18 0 0 8320 0 6 30 0 0 3
177 1451
177 1455
306 1455
0 2 19 0 0 8192 0 0 32 23 0 4
286 1359
294 1359
294 1397
304 1397
1 1 19 0 0 8192 0 7 32 0 0 5
174 1327
174 1359
286 1359
286 1379
304 1379
1 2 18 0 0 0 0 6 31 0 0 4
177 1451
188 1451
188 1323
302 1323
1 1 19 0 0 8320 0 7 31 0 0 3
174 1327
174 1305
302 1305
3 0 20 0 0 0 0 33 0 0 28 2
1009 1020
1009 1020
3 0 21 0 0 0 0 34 0 0 33 2
436 989
436 989
0 1 20 0 0 4224 0 0 35 0 0 3
1006 1020
1058 1020
1058 1016
1 2 22 0 0 4224 0 8 33 0 0 4
880 1078
949 1078
949 1029
954 1029
1 1 23 0 0 4224 0 9 33 0 0 4
872 958
949 958
949 1011
954 1011
4 1 24 0 0 4224 0 37 36 0 0 3
566 989
614 989
614 980
3 3 25 0 0 4224 0 38 37 0 0 4
296 1037
509 1037
509 998
520 998
0 2 21 0 0 4224 0 0 37 0 0 2
433 989
521 989
3 1 26 0 0 4224 0 39 37 0 0 4
294 904
509 904
509 980
520 980
1 2 27 0 0 4224 0 10 34 0 0 4
162 1119
371 1119
371 998
381 998
1 1 28 0 0 4224 0 12 34 0 0 2
151 980
381 980
1 2 29 0 0 4224 0 13 39 0 0 2
148 913
249 913
1 1 29 0 0 0 0 13 41 0 0 4
148 913
198 913
198 895
204 895
1 2 30 0 0 4224 0 11 38 0 0 2
155 1046
251 1046
1 1 30 0 0 0 0 11 40 0 0 4
155 1046
201 1046
201 1028
205 1028
1 2 31 0 0 4224 0 38 40 0 0 2
251 1028
241 1028
1 2 32 0 0 4224 0 39 41 0 0 2
249 895
240 895
3 1 33 0 0 4224 0 43 42 0 0 3
693 721
743 721
743 713
1 2 34 0 0 4224 0 14 44 0 0 2
154 784
265 784
3 2 35 0 0 4224 0 44 43 0 0 4
316 775
634 775
634 730
642 730
3 1 36 0 0 4224 0 45 43 0 0 4
477 680
634 680
634 712
642 712
0 1 37 0 0 4224 0 0 44 51 0 3
181 586
181 766
265 766
3 1 38 0 0 4224 0 46 45 0 0 4
315 595
418 595
418 671
426 671
1 2 39 0 0 4224 0 15 45 0 0 4
154 676
418 676
418 689
426 689
0 2 37 0 0 0 0 0 46 51 0 3
217 586
217 604
264 604
1 1 37 0 0 0 0 16 46 0 0 2
151 586
264 586
2 1 40 0 0 4224 0 49 47 0 0 5
518 479
609 479
609 486
621 486
621 478
1 1 41 0 0 4096 0 49 17 0 0 4
482 479
173 479
173 281
154 281
2 1 42 0 0 4224 0 50 48 0 0 5
516 415
606 415
606 421
618 421
618 413
1 1 43 0 0 4096 0 18 50 0 0 4
149 144
455 144
455 415
480 415
3 1 44 0 0 4224 0 57 51 0 0 5
525 347
602 347
602 364
614 364
614 356
3 1 45 0 0 4224 0 58 52 0 0 5
525 277
594 277
594 294
606 294
606 286
3 1 46 0 0 4224 0 59 53 0 0 5
525 214
588 214
588 233
600 233
600 225
3 1 47 0 0 4224 0 60 54 0 0 5
519 162
586 162
586 174
598 174
598 166
3 1 48 0 0 4224 0 61 55 0 0 5
521 106
581 106
581 120
593 120
593 112
1 2 41 0 0 0 0 17 57 0 0 4
154 281
185 281
185 356
470 356
1 1 43 0 0 12288 0 18 57 0 0 4
149 144
161 144
161 338
470 338
1 1 43 0 0 4096 0 18 58 0 0 4
149 144
468 144
468 268
476 268
1 2 41 0 0 8320 0 17 58 0 0 5
154 281
154 287
468 287
468 286
476 286
1 2 41 0 0 0 0 17 59 0 0 4
154 281
170 281
170 223
473 223
0 1 43 0 0 0 0 0 59 68 0 3
289 144
289 205
473 205
1 2 41 0 0 0 0 17 61 0 0 4
154 281
246 281
246 115
470 115
0 1 43 0 0 0 0 0 61 70 0 4
149 144
462 144
462 97
470 97
1 2 41 0 0 0 0 17 60 0 0 4
154 281
465 281
465 171
473 171
0 1 43 0 0 8320 0 0 60 72 0 4
149 144
149 154
473 154
473 153
3 1 49 0 0 4224 0 62 56 0 0 3
514 45
592 45
592 37
1 1 43 0 0 0 0 62 18 0 0 4
469 36
171 36
171 144
149 144
2 1 41 0 0 0 0 62 17 0 0 4
469 54
183 54
183 281
154 281
32
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
94 266 123 290
104 274 112 290
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
97 126 122 150
105 134 113 150
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 91
924 42 1097 186
934 50 1086 162
91 Tabela Verdade AND:

A    B    Sa�da:
0    0    0
0    1    0
1    0    0
1    1    1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 92
929 195 1110 339
939 203 1099 315
92 Tabela Verdade NAND:

A    B    Sa�da:
0    0    1
0    1    1
1    0    1
1    1    0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 90
920 364 1085 508
930 372 1074 484
90 Tabela Verdade OR:

A    B    Sa�da:
0    0    0
0    1    1
1    0    1
1    1    1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 91
1144 43 1317 187
1154 51 1306 163
91 Tabela Verdade NOR:

A    B    Sa�da:
0    0    1
0    1    0
1    0    0
1    1    0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 91
1144 193 1317 337
1154 201 1306 313
91 Tabela Verdade XOR:

A    B    Sa�da:
0    0    0
0    1    1
1    0    1
1    1    0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 92
1147 362 1328 506
1157 370 1317 482
92 Tabela Verdade NXOR:

A    B    Sa�da:
0    0    1
0    1    0
1    0    0
1    1    1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 88
711 44 916 148
721 52 905 132
88 Tabela Verdade NOT:

A    Sa�da   B    Sa�da
0    1       0    1
1    0       1    0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
63 10 140 34
73 18 129 34
7 a) e b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
90 892 119 916
100 900 108 916
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
93 955 122 979
103 963 111 979
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
96 1017 125 1041
106 1025 114 1041
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
104 1104 133 1128
114 1112 122 1128
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
719 983 748 1007
729 991 737 1007
1 =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
815 941 844 965
825 949 833 965
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
824 1061 853 1085
834 1069 842 1085
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 42
75 820 432 844
85 828 421 844
42 c.1,1)Simplificando: m(0,2,5,7,8,10,13,15)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
82 570 111 594
92 578 100 594
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
86 760 115 784
96 768 104 784
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
88 660 117 684
98 668 106 684
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 51
100 1225 529 1249
110 1233 518 1249
51 c.2,1) Aplicando somente portas NAND no 1� Circuito
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
109 1311 138 1335
119 1319 127 1335
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
112 1437 141 1461
122 1445 130 1461
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 51
35 503 464 527
45 511 453 527
51 c.2,1) Aplicando somente portas NAND no 2� Circuito
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 33
124 1570 409 1594
134 1578 398 1594
33 C.1,2)Simplificando o 2� Circuito
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
143 1659 172 1683
153 1667 161 1683
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
144 1725 173 1749
154 1733 162 1749
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
142 1781 171 1805
152 1789 160 1805
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
93 1890 130 1914
103 1898 119 1914
2 d)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
215 1895 244 1919
225 1903 233 1919
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
218 2028 247 2052
228 2036 236 2052
1 B
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
