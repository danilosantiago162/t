CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 50 30 100 10
176 80 1364 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499192 0.500000
176 80 1364 388
9437202 0
0
6 Title:
5 Name:
0
0
0
43
13 Logic Switch~
5 171 298 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45417.6 0
0
13 Logic Switch~
5 168 230 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45417.6 0
0
13 Logic Switch~
5 172 170 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
45417.6 0
0
13 Logic Switch~
5 173 112 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
45417.6 0
0
14 Logic Display~
6 888 82 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
45417.6 0
0
14 Logic Display~
6 898 643 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
45417.6 0
0
14 Logic Display~
6 897 587 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
45417.6 0
0
14 Logic Display~
6 898 523 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
45417.6 0
0
14 Logic Display~
6 894 471 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
45417.6 0
0
14 Logic Display~
6 891 403 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
45417.6 0
0
14 Logic Display~
6 888 345 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
45417.6 0
0
14 Logic Display~
6 887 263 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
45417.6 0
0
14 Logic Display~
6 887 207 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
45417.6 0
0
14 Logic Display~
6 887 150 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4597 0 0
2
45417.6 0
0
5 4049~
219 406 289 0 2 22
0 22 12
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 9 0
1 U
3835 0 0
2
45417.6 0
0
5 4049~
219 396 546 0 2 22
0 22 13
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 9 0
1 U
3670 0 0
2
45417.6 0
0
5 4049~
219 396 493 0 2 22
0 22 14
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 9 0
1 U
5616 0 0
2
45417.6 0
0
5 4049~
219 405 230 0 2 22
0 22 15
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 8 0
1 U
9323 0 0
2
45417.6 0
0
5 4049~
219 498 677 0 2 22
0 21 16
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 8 0
1 U
317 0 0
2
45417.6 0
0
5 4049~
219 496 555 0 2 22
0 21 17
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 8 0
1 U
3108 0 0
2
45417.6 0
0
5 4049~
219 489 435 0 2 22
0 21 18
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 8 0
1 U
4299 0 0
2
45417.6 0
0
5 4049~
219 484 298 0 2 22
0 21 19
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 8 0
1 U
9672 0 0
2
45417.6 0
0
5 4049~
219 487 181 0 2 22
0 21 20
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 8 0
1 U
7876 0 0
2
45417.6 0
0
5 4049~
219 713 650 0 2 22
0 33 23
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 7 0
1 U
6369 0 0
2
45417.6 0
0
5 4049~
219 709 593 0 2 22
0 33 24
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 7 0
1 U
9172 0 0
2
45417.6 0
0
5 4049~
219 317 537 0 2 22
0 25 28
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 7 0
1 U
7100 0 0
2
45417.6 0
0
5 4049~
219 314 484 0 2 22
0 25 29
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 7 0
1 U
3820 0 0
2
45417.6 0
0
5 4049~
219 315 417 0 2 22
0 25 30
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 7 0
1 U
7678 0 0
2
45417.6 0
0
5 4049~
219 316 360 0 2 22
0 25 31
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 6 0
1 U
961 0 0
2
45417.6 0
0
5 4049~
219 214 298 0 2 22
0 26 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 6 0
1 U
3178 0 0
2
45417.6 0
0
5 4049~
219 215 230 0 2 22
0 27 22
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 6 0
1 U
3409 0 0
2
45417.6 0
0
5 4049~
219 215 170 0 2 22
0 32 25
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 6 0
1 U
3951 0 0
2
45417.6 0
0
5 4049~
219 217 112 0 2 22
0 34 33
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 6 0
1 U
8885 0 0
2
45417.6 0
0
5 4082~
219 855 663 0 5 22
0 23 25 22 16 11
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
3780 0 0
2
45417.6 0
0
5 4082~
219 855 606 0 5 22
0 24 25 22 21 10
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
9265 0 0
2
45417.6 0
0
5 4082~
219 854 541 0 5 22
0 33 28 13 17 9
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
9442 0 0
2
45417.6 0
0
5 4082~
219 854 488 0 5 22
0 33 29 14 21 8
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
9424 0 0
2
45417.6 0
0
5 4082~
219 852 421 0 5 22
0 33 30 22 18 7
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
9968 0 0
2
45417.6 0
0
5 4082~
219 853 364 0 5 22
0 33 31 22 21 6
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
9281 0 0
2
45417.6 0
0
5 4082~
219 851 284 0 5 22
0 33 25 12 19 5
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
8464 0 0
2
45417.6 0
0
5 4082~
219 850 225 0 5 22
0 33 25 15 21 4
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
7168 0 0
2
45417.6 0
0
5 4082~
219 850 167 0 5 22
0 33 25 22 20 3
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
3171 0 0
2
45417.6 0
0
5 4082~
219 849 101 0 5 22
0 33 25 22 21 2
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
4139 0 0
2
45417.6 0
0
69
5 1 2 0 0 4240 0 43 5 0 0 3
870 101
888 101
888 100
5 1 3 0 0 4224 0 42 14 0 0 3
871 167
887 167
887 168
5 1 4 0 0 4224 0 41 13 0 0 2
871 225
887 225
5 1 5 0 0 4224 0 40 12 0 0 3
872 284
887 284
887 281
5 1 6 0 0 4224 0 39 11 0 0 3
874 364
888 364
888 363
5 1 7 0 0 4224 0 38 10 0 0 2
873 421
891 421
5 1 8 0 0 4224 0 37 9 0 0 3
875 488
894 488
894 489
5 1 9 0 0 4224 0 36 8 0 0 2
875 541
898 541
5 1 10 0 0 4224 0 35 7 0 0 3
876 606
897 606
897 605
5 1 11 0 0 4224 0 34 6 0 0 3
876 663
898 663
898 661
2 3 12 0 0 4224 0 15 40 0 0 2
427 289
827 289
2 3 13 0 0 4224 0 16 36 0 0 2
417 546
830 546
2 3 14 0 0 4224 0 17 37 0 0 2
417 493
830 493
2 3 15 0 0 4224 0 18 41 0 0 2
426 230
826 230
2 4 16 0 0 4224 0 19 34 0 0 2
519 677
831 677
2 4 17 0 0 4224 0 20 36 0 0 2
517 555
830 555
2 4 18 0 0 4224 0 21 38 0 0 2
510 435
828 435
2 4 19 0 0 4224 0 22 40 0 0 2
505 298
827 298
2 4 20 0 0 4224 0 23 42 0 0 2
508 181
826 181
0 4 21 0 0 8192 0 0 43 29 0 3
452 183
452 115
825 115
4 0 21 0 0 4096 0 41 0 0 29 2
826 239
452 239
0 1 21 0 0 0 0 0 22 29 0 2
452 298
469 298
4 0 21 0 0 4096 0 39 0 0 28 2
829 378
452 378
0 1 21 0 0 0 0 0 21 28 0 2
452 435
474 435
4 0 21 0 0 4096 0 37 0 0 28 2
830 502
452 502
0 1 21 0 0 0 0 0 20 28 0 2
452 555
481 555
4 0 21 0 0 4224 0 35 0 0 28 2
831 620
452 620
0 1 21 0 0 0 0 0 19 29 0 3
452 298
452 677
483 677
2 1 21 0 0 0 0 30 23 0 0 6
235 298
452 298
452 305
452 305
452 181
472 181
3 0 22 0 0 4096 0 42 0 0 41 2
826 172
353 172
0 1 22 0 0 0 0 0 18 41 0 2
353 230
390 230
0 1 22 0 0 0 0 0 15 40 0 4
353 290
358 290
358 289
391 289
3 0 22 0 0 4096 0 39 0 0 40 2
829 369
353 369
3 0 22 0 0 0 0 38 0 0 40 2
828 426
353 426
0 1 22 0 0 0 0 0 17 40 0 4
353 494
358 494
358 493
381 493
0 1 22 0 0 0 0 0 16 40 0 2
353 546
381 546
3 0 22 0 0 4224 0 35 0 0 40 2
831 611
353 611
2 1 23 0 0 4224 0 24 34 0 0 2
734 650
831 650
2 1 24 0 0 4224 0 25 35 0 0 2
730 593
831 593
0 3 22 0 0 0 0 0 34 41 0 3
353 230
353 668
831 668
2 3 22 0 0 0 0 31 43 0 0 4
236 230
353 230
353 106
825 106
2 0 25 0 0 4224 0 35 0 0 56 2
831 602
286 602
1 1 26 0 0 4224 0 1 30 0 0 2
183 298
199 298
1 1 27 0 0 4224 0 2 31 0 0 2
180 230
200 230
2 2 28 0 0 4224 0 26 36 0 0 2
338 537
830 537
0 1 25 0 0 0 0 0 26 56 0 2
286 537
302 537
2 2 29 0 0 4224 0 27 37 0 0 2
335 484
830 484
1 0 25 0 0 0 0 27 0 0 56 2
299 484
286 484
2 2 30 0 0 4224 0 28 38 0 0 2
336 417
828 417
1 0 25 0 0 0 0 28 0 0 56 2
300 417
286 417
2 2 31 0 0 4224 0 29 39 0 0 2
337 360
829 360
1 0 25 0 0 0 0 29 0 0 56 2
301 360
286 360
2 0 25 0 0 0 0 40 0 0 56 2
827 280
286 280
2 0 25 0 0 0 0 41 0 0 56 2
826 221
286 221
2 0 25 0 0 0 0 42 0 0 57 2
826 163
286 163
0 2 25 0 0 0 0 0 34 57 0 3
286 170
286 659
831 659
2 2 25 0 0 0 0 32 43 0 0 4
236 170
286 170
286 97
825 97
1 1 32 0 0 4224 0 3 32 0 0 2
184 170
200 170
0 1 33 0 0 4096 0 0 38 63 0 2
267 408
828 408
0 1 33 0 0 4224 0 0 37 63 0 2
267 475
830 475
0 1 33 0 0 0 0 0 36 63 0 2
267 528
830 528
0 1 33 0 0 0 0 0 25 63 0 2
267 593
694 593
0 1 33 0 0 0 0 0 24 64 0 3
267 351
267 650
698 650
0 1 33 0 0 0 0 0 39 65 0 3
267 271
267 351
829 351
0 1 33 0 0 0 0 0 40 66 0 3
267 212
267 271
827 271
0 1 33 0 0 0 0 0 41 67 0 3
267 154
267 212
826 212
0 1 33 0 0 0 0 0 42 68 0 3
267 112
267 154
826 154
2 1 33 0 0 0 0 33 43 0 0 4
238 112
267 112
267 88
825 88
1 1 34 0 0 4224 0 4 33 0 0 2
185 112
202 112
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
123 277 148 301
131 285 139 301
1 Z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
122 225 147 249
130 233 138 249
1 W
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
122 151 147 175
130 159 138 175
1 Y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
120 95 145 119
128 103 136 119
1 X
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
