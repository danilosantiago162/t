CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 90 30 100 10
176 80 1364 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 37 302 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
523 0 0
2
45423.8 0
0
13 Logic Switch~
5 42 245 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-3 -27 4 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6748 0 0
2
45423.8 0
0
13 Logic Switch~
5 39 190 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -17 8 -9
1 B
-3 -25 4 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6901 0 0
2
45423.8 0
0
13 Logic Switch~
5 36 129 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
842 0 0
2
45423.8 0
0
8 4-In OR~
219 402 439 0 5 22
0 16 20 9 2 19
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
3277 0 0
2
45423.9 0
0
8 2-In OR~
219 240 633 0 3 22
0 6 3 4
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U2D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
4212 0 0
2
45423.9 0
0
9 2-In AND~
219 337 605 0 3 22
0 5 4 2
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
4720 0 0
2
45423.9 0
0
9 2-In AND~
219 271 586 0 3 22
0 8 7 5
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
5551 0 0
2
45423.9 0
0
5 4049~
219 98 245 0 2 22
0 15 7
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 4 0
1 U
6986 0 0
2
45423.8 0
0
8 2-In OR~
219 229 381 0 3 22
0 8 7 17
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U2C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8745 0 0
2
45423.8 0
0
5 4049~
219 86 129 0 2 22
0 13 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 4 0
1 U
9592 0 0
2
45423.8 0
0
9 2-In AND~
219 298 372 0 3 22
0 18 17 16
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
8748 0 0
2
45423.8 0
0
9 2-In AND~
219 124 458 0 3 22
0 13 12 21
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
7168 0 0
2
45423.8 0
0
9 2-In AND~
219 236 346 0 3 22
0 6 3 18
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
631 0 0
2
45423.8 0
0
9 2-In AND~
219 178 529 0 3 22
0 11 10 9
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9466 0 0
2
45423.8 0
0
5 4030~
219 117 414 0 3 22
0 15 14 22
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
3266 0 0
2
45423.8 0
0
5 4030~
219 115 507 0 3 22
0 13 12 11
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
7693 0 0
2
45423.8 0
0
9 2-In AND~
219 121 554 0 3 22
0 15 14 10
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3723 0 0
2
45423.8 0
0
9 2-In AND~
219 186 437 0 3 22
0 22 21 20
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3440 0 0
2
45423.8 0
0
5 4049~
219 104 302 0 2 22
0 14 3
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 4 0
1 U
6263 0 0
2
45423.8 0
0
5 4049~
219 93 164 0 2 22
0 12 6
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 4 0
1 U
4900 0 0
2
45423.8 0
0
8 3-In OR~
219 460 220 0 4 22
0 24 26 25 23
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
8783 0 0
2
45423.8 0
0
8 2-In OR~
219 165 274 0 3 22
0 7 3 28
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3221 0 0
2
45423.8 0
0
8 2-In OR~
219 170 164 0 3 22
0 8 6 27
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3215 0 0
2
45423.8 0
0
9 2-In AND~
219 324 149 0 3 22
0 8 6 24
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7903 0 0
2
45423.8 0
0
9 2-In AND~
219 266 220 0 3 22
0 27 28 26
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7121 0 0
2
45423.8 0
0
9 2-In AND~
219 325 270 0 3 22
0 7 3 25
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4484 0 0
2
45423.8 0
0
14 Logic Display~
6 646 136 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5996 0 0
2
45423.8 0
0
14 Logic Display~
6 536 137 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7804 0 0
2
45423.8 0
0
47
4 3 2 0 0 8320 0 5 7 0 0 4
385 453
366 453
366 605
358 605
0 2 3 0 0 4240 0 0 6 21 0 3
149 355
149 642
227 642
2 3 4 0 0 12416 0 7 6 0 0 4
313 614
309 614
309 633
273 633
3 1 5 0 0 4224 0 8 7 0 0 4
292 586
305 586
305 596
313 596
0 1 6 0 0 4224 0 0 6 22 0 3
125 337
125 624
227 624
0 2 7 0 0 8320 0 0 8 19 0 4
132 381
144 381
144 595
247 595
0 1 8 0 0 8192 0 0 8 20 0 4
120 372
155 372
155 577
247 577
0 1 7 0 0 0 0 0 23 47 0 5
141 245
141 249
144 249
144 265
152 265
3 3 9 0 0 4224 0 15 5 0 0 5
199 529
359 529
359 445
385 445
385 444
3 2 10 0 0 8320 0 18 15 0 0 4
142 554
146 554
146 538
154 538
3 1 11 0 0 4224 0 17 15 0 0 3
148 507
148 520
154 520
0 2 12 0 0 4096 0 0 17 29 0 3
71 466
71 516
99 516
0 1 13 0 0 4096 0 0 17 30 0 3
66 447
66 498
99 498
0 2 14 0 0 4224 0 0 18 27 0 3
84 423
84 563
97 563
0 1 15 0 0 4096 0 0 18 28 0 3
78 405
78 545
97 545
3 1 16 0 0 8320 0 12 5 0 0 5
319 372
359 372
359 427
385 427
385 426
3 2 17 0 0 4224 0 10 12 0 0 2
262 381
274 381
3 1 18 0 0 8320 0 14 12 0 0 4
257 346
266 346
266 363
274 363
0 2 7 0 0 0 0 0 10 47 0 5
132 245
132 243
132 243
132 390
216 390
0 1 8 0 0 4224 0 0 10 38 0 3
120 129
120 372
216 372
0 2 3 0 0 0 0 0 14 33 0 3
129 302
129 355
212 355
0 1 6 0 0 0 0 0 14 37 0 3
125 189
125 337
212 337
5 1 19 0 0 12416 0 5 28 0 0 4
435 439
435 438
646 438
646 154
3 2 20 0 0 4224 0 19 5 0 0 5
207 437
359 437
359 436
385 436
385 435
3 2 21 0 0 8320 0 13 19 0 0 4
145 458
154 458
154 446
162 446
3 1 22 0 0 8320 0 16 19 0 0 4
150 414
154 414
154 428
162 428
0 2 14 0 0 0 0 0 16 34 0 3
84 302
84 423
101 423
0 1 15 0 0 4224 0 0 16 35 0 3
78 245
78 405
101 405
0 2 12 0 0 4224 0 0 13 36 0 3
71 190
71 467
100 467
0 1 13 0 0 4224 0 0 13 31 0 3
66 129
66 449
100 449
1 1 13 0 0 128 0 11 4 0 0 2
71 129
48 129
0 2 3 0 0 128 0 0 27 33 0 4
144 302
293 302
293 279
301 279
2 2 3 0 0 0 0 20 23 0 0 4
125 302
144 302
144 283
152 283
1 1 14 0 0 0 0 20 1 0 0 2
89 302
49 302
1 1 15 0 0 128 0 2 9 0 0 2
54 245
83 245
1 1 12 0 0 128 0 3 21 0 0 4
51 190
71 190
71 164
78 164
2 2 6 0 0 0 0 21 24 0 0 8
114 164
125 164
125 189
138 189
138 190
138 190
138 173
157 173
2 1 8 0 0 0 0 11 24 0 0 6
107 129
179 129
179 129
138 129
138 155
157 155
4 1 23 0 0 8320 0 22 29 0 0 3
493 220
536 220
536 155
3 1 24 0 0 8320 0 25 22 0 0 4
345 149
390 149
390 211
447 211
0 1 8 0 0 128 0 0 25 38 0 4
179 129
209 129
209 140
300 140
0 2 6 0 0 128 0 0 25 37 0 4
138 190
292 190
292 158
300 158
3 3 25 0 0 12416 0 27 22 0 0 4
346 270
390 270
390 229
447 229
3 2 26 0 0 4224 0 26 22 0 0 2
287 220
448 220
3 1 27 0 0 8320 0 24 26 0 0 4
203 164
226 164
226 211
242 211
3 2 28 0 0 8320 0 23 26 0 0 4
198 274
226 274
226 229
242 229
2 1 7 0 0 128 0 9 27 0 0 4
119 245
293 245
293 261
301 261
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
