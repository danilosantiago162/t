CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 485
9437202 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 65 255 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8745 0 0
2
45435.7 0
0
13 Logic Switch~
5 63 322 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9592 0 0
2
45435.7 0
0
13 Logic Switch~
5 55 394 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8748 0 0
2
45435.7 0
0
13 Logic Switch~
5 56 465 0 1 11
0 31
0
0 0 21360 0
2 0V
-7 -16 7 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7168 0 0
2
45435.7 0
0
13 Logic Switch~
5 49 55 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
631 0 0
2
45435.7 0
0
13 Logic Switch~
5 74 55 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9466 0 0
2
45435.7 0
0
13 Logic Switch~
5 101 55 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3266 0 0
2
45435.7 0
0
13 Logic Switch~
5 123 56 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7693 0 0
2
45435.7 0
0
8 2-In OR~
219 693 274 0 3 22
0 10 9 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3723 0 0
2
45435.7 0
0
8 2-In OR~
219 690 206 0 3 22
0 15 14 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3440 0 0
2
45435.7 0
0
5 7405~
219 527 169 0 2 22
0 5 12
0
0 0 624 0
6 74LS05
-21 -24 21 -16
3 U8C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 6 0
65 0 0 0 6 3 6 0
1 U
6263 0 0
2
45435.7 0
0
5 7405~
219 556 333 0 2 22
0 2 7
0
0 0 624 0
6 74LS05
-21 -24 21 -16
3 U8B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 6 0
65 0 0 0 6 2 6 0
1 U
4900 0 0
2
45435.7 0
0
5 7405~
219 554 215 0 2 22
0 11 6
0
0 0 624 0
6 74LS05
-21 -24 21 -16
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 6 0
65 0 0 0 6 1 6 0
1 U
8783 0 0
2
45435.7 0
0
9 2-In AND~
219 645 264 0 3 22
0 12 2 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3221 0 0
2
45435.7 0
0
9 2-In AND~
219 646 225 0 3 22
0 12 11 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3215 0 0
2
45435.7 0
0
9 2-In AND~
219 645 295 0 3 22
0 2 11 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
7903 0 0
2
45435.7 0
0
5 7415~
219 614 324 0 4 22
0 5 6 7 4
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 4 0
1 U
7121 0 0
2
45435.7 0
0
5 7415~
219 654 193 0 4 22
0 5 2 6 15
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 4 0
1 U
4484 0 0
2
45435.7 0
0
8 2-In OR~
219 912 112 0 3 22
0 19 18 17
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5996 0 0
2
45435.7 0
0
9 2-In AND~
219 852 137 0 3 22
0 21 20 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7804 0 0
2
45435.7 0
0
9 2-In AND~
219 851 91 0 3 22
0 21 22 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5523 0 0
2
45435.7 0
0
12 Hex Display~
7 670 360 0 18 19
10 17 35 36 37 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
3330 0 0
2
45435.7 0
0
12 Hex Display~
7 716 361 0 18 19
10 16 13 8 4 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3465 0 0
2
45435.7 0
0
6 74LS83
105 709 116 0 14 29
0 30 29 28 27 26 25 24 23 38
21 22 20 39 3
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
8396 0 0
2
45435.7 0
0
9 2-In XOR~
219 189 474 0 3 22
0 31 3 23
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3685 0 0
2
45435.7 0
0
9 2-In XOR~
219 193 403 0 3 22
0 32 3 24
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7849 0 0
2
45435.7 0
0
9 2-In XOR~
219 186 331 0 3 22
0 33 3 25
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6343 0 0
2
45435.7 0
0
9 2-In XOR~
219 183 264 0 3 22
0 34 3 26
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7376 0 0
2
45435.7 0
0
6 74LS83
105 462 206 0 14 29
0 30 29 28 27 26 25 24 23 40
5 2 11 16 3
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
9156 0 0
2
45435.7 5
0
55
0 1 2 0 0 4112 0 0 16 22 0 3
614 192
614 286
621 286
14 0 3 0 0 8192 0 24 0 0 43 4
741 161
741 248
495 248
495 251
4 4 4 0 0 8320 0 17 23 0 0 6
635 324
635 317
764 317
764 404
707 404
707 385
1 10 5 0 0 8192 0 17 29 0 0 4
590 315
505 315
505 197
494 197
0 2 6 0 0 4224 0 0 17 20 0 3
583 215
583 324
590 324
0 1 2 0 0 4224 0 0 12 22 0 3
511 206
511 333
541 333
3 2 7 0 0 4224 0 17 12 0 0 2
590 333
577 333
3 3 8 0 0 8320 0 9 23 0 0 5
726 274
743 274
743 398
713 398
713 385
3 2 9 0 0 8320 0 16 9 0 0 4
666 295
672 295
672 283
680 283
3 1 10 0 0 12416 0 14 9 0 0 4
666 264
672 264
672 265
680 265
0 2 11 0 0 4096 0 0 16 17 0 3
562 234
562 304
621 304
0 2 2 0 0 0 0 0 14 22 0 3
589 192
589 273
621 273
0 1 12 0 0 4224 0 0 14 15 0 3
600 169
600 255
621 255
3 2 13 0 0 8320 0 10 23 0 0 5
723 206
738 206
738 393
719 393
719 385
2 1 12 0 0 0 0 11 15 0 0 4
548 169
609 169
609 216
622 216
0 1 5 0 0 0 0 0 11 23 0 3
495 197
495 169
512 169
0 2 11 0 0 8320 0 0 15 21 0 3
530 215
530 234
622 234
3 2 14 0 0 4224 0 15 10 0 0 3
667 225
667 215
677 215
4 1 15 0 0 8320 0 18 10 0 0 4
675 193
676 193
676 197
677 197
2 3 6 0 0 0 0 13 18 0 0 4
575 215
583 215
583 202
630 202
12 1 11 0 0 0 0 29 13 0 0 2
494 215
539 215
11 2 2 0 0 0 0 29 18 0 0 5
494 206
540 206
540 192
630 192
630 193
10 1 5 0 0 4224 0 29 18 0 0 4
494 197
619 197
619 184
630 184
13 1 16 0 0 12416 0 29 23 0 0 5
494 224
525 224
525 413
725 413
725 385
3 1 17 0 0 8320 0 19 22 0 0 5
945 112
949 112
949 422
679 422
679 384
3 2 18 0 0 4224 0 20 19 0 0 4
873 137
891 137
891 121
899 121
3 1 19 0 0 4224 0 21 19 0 0 4
872 91
891 91
891 103
899 103
12 2 20 0 0 4224 0 24 20 0 0 4
741 125
820 125
820 146
828 146
0 1 21 0 0 8192 0 0 20 31 0 3
769 107
769 128
828 128
11 2 22 0 0 4224 0 24 21 0 0 4
741 116
814 116
814 100
827 100
10 1 21 0 0 4224 0 24 21 0 0 4
741 107
819 107
819 82
827 82
0 8 23 0 0 4224 0 0 24 48 0 3
361 474
361 143
677 143
0 7 24 0 0 8320 0 0 24 49 0 3
369 403
369 134
677 134
0 6 25 0 0 8320 0 0 24 50 0 3
378 331
378 125
677 125
0 5 26 0 0 8320 0 0 24 51 0 3
387 264
387 116
677 116
4 0 27 0 0 4224 0 24 0 0 55 2
677 107
123 107
3 0 28 0 0 4224 0 24 0 0 54 2
677 98
101 98
2 0 29 0 0 4224 0 24 0 0 53 2
677 89
74 89
1 0 30 0 0 4224 0 24 0 0 52 2
677 80
49 80
0 2 3 0 0 4224 0 0 28 43 0 4
495 289
153 289
153 273
167 273
0 2 3 0 0 0 0 0 27 43 0 4
495 357
155 357
155 340
170 340
0 2 3 0 0 0 0 0 26 43 0 4
495 428
159 428
159 412
177 412
14 2 3 0 0 0 0 29 25 0 0 6
494 251
495 251
495 501
165 501
165 483
173 483
1 1 31 0 0 4224 0 4 25 0 0 2
68 465
173 465
1 1 32 0 0 4224 0 3 26 0 0 2
67 394
177 394
1 1 33 0 0 4224 0 2 27 0 0 2
75 322
170 322
1 1 34 0 0 4224 0 1 28 0 0 2
77 255
167 255
3 8 23 0 0 0 0 25 29 0 0 4
222 474
404 474
404 233
430 233
3 7 24 0 0 0 0 26 29 0 0 4
226 403
409 403
409 224
430 224
3 6 25 0 0 0 0 27 29 0 0 4
219 331
414 331
414 215
430 215
3 5 26 0 0 0 0 28 29 0 0 4
216 264
419 264
419 206
430 206
1 1 30 0 0 0 0 5 29 0 0 3
49 67
49 170
430 170
1 2 29 0 0 0 0 6 29 0 0 3
74 67
74 179
430 179
1 3 28 0 0 0 0 7 29 0 0 3
101 67
101 188
430 188
1 4 27 0 0 0 0 8 29 0 0 3
123 68
123 197
430 197
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
