CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1364 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
38
13 Logic Switch~
5 132 618 0 1 11
0 7
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45435.7 7
0
13 Logic Switch~
5 365 601 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45435.7 6
0
13 Logic Switch~
5 388 601 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
45435.7 5
0
13 Logic Switch~
5 157 619 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
45435.7 4
0
13 Logic Switch~
5 181 616 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
45435.7 3
0
13 Logic Switch~
5 411 601 0 1 11
0 5
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B1
-4 -32 10 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
45435.7 2
0
13 Logic Switch~
5 203 615 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
45435.7 1
0
13 Logic Switch~
5 433 601 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 B0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
45435.7 0
0
9 2-In AND~
219 185 749 0 3 22
0 7 38 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
4747 0 0
2
45435.7 37
0
5 4049~
219 123 758 0 2 22
0 8 38
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 14 0
1 U
972 0 0
2
45435.7 36
0
9 2-In AND~
219 190 798 0 3 22
0 8 37 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3472 0 0
2
45435.7 35
0
5 4049~
219 125 725 0 2 22
0 7 37
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 14 0
1 U
9998 0 0
2
45435.7 34
0
5 4049~
219 357 688 0 2 22
0 10 36
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 14 0
1 U
3536 0 0
2
45435.7 33
0
5 7415~
219 453 774 0 4 22
0 36 31 9 35
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U15C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 13 0
1 U
4597 0 0
2
45435.7 32
0
8 2-In OR~
219 496 807 0 3 22
0 35 33 25
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U14D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
3835 0 0
2
45435.7 31
0
5 7415~
219 458 717 0 4 22
0 10 34 32 30
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U15B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 13 0
1 U
3670 0 0
2
45435.7 30
0
5 4049~
219 363 743 0 2 22
0 9 34
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16C
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 14 0
1 U
5616 0 0
2
45435.7 29
0
5 4049~
219 264 799 0 2 22
0 33 32
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 14 0
1 U
9323 0 0
2
45435.7 28
0
5 4049~
219 287 770 0 2 22
0 29 31
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 14 0
1 U
317 0 0
2
45435.7 27
0
8 2-In OR~
219 517 726 0 3 22
0 30 29 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U14C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
3108 0 0
2
45435.7 26
0
8 2-In OR~
219 884 722 0 3 22
0 22 21 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U14B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
4299 0 0
2
45435.7 25
0
5 4049~
219 613 770 0 2 22
0 21 23
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U13F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 11 0
1 U
9672 0 0
2
45435.7 24
0
5 4049~
219 572 787 0 2 22
0 25 24
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U13E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 11 0
1 U
7876 0 0
2
45435.7 23
0
5 4049~
219 740 720 0 2 22
0 5 26
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U13D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 11 0
1 U
6369 0 0
2
45435.7 22
0
5 7415~
219 805 678 0 4 22
0 6 26 24 22
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U15A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 13 0
1 U
9172 0 0
2
45435.7 21
0
8 2-In OR~
219 796 811 0 3 22
0 27 25 17
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U14A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
7100 0 0
2
45435.7 20
0
5 7415~
219 750 770 0 4 22
0 28 23 5 27
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U12C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 10 0
1 U
3820 0 0
2
45435.7 19
0
5 4049~
219 589 695 0 2 22
0 6 28
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U13C
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 11 0
1 U
7678 0 0
2
45435.7 18
0
8 2-In OR~
219 1092 734 0 3 22
0 14 13 12
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
961 0 0
2
45435.7 17
0
5 4049~
219 958 777 0 2 22
0 13 15
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U13B
-13 -17 15 -9
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 11 0
1 U
3178 0 0
2
45435.7 16
0
5 4049~
219 861 788 0 2 22
0 17 16
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U13A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 11 0
1 U
3409 0 0
2
45435.7 15
0
5 4049~
219 970 722 0 2 22
0 4 18
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 9 0
1 U
3951 0 0
2
45435.7 14
0
5 7415~
219 1046 702 0 4 22
0 3 18 16 14
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U12B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 10 0
1 U
8885 0 0
2
45435.7 13
0
8 2-In OR~
219 1092 786 0 3 22
0 19 17 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3780 0 0
2
45435.7 12
0
5 7415~
219 1039 777 0 4 22
0 20 15 4 19
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U12A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 10 0
1 U
9265 0 0
2
45435.7 11
0
5 4049~
219 970 674 0 2 22
0 3 20
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 9 0
1 U
9442 0 0
2
45435.7 10
0
14 Logic Display~
6 1137 592 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 X
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9424 0 0
2
45435.7 9
0
14 Logic Display~
6 1169 592 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9968 0 0
2
45435.7 8
0
50
1 1 3 0 0 8320 0 7 33 0 0 7
203 627
203 635
950 635
950 694
950 694
950 693
1022 693
1 1 4 0 0 8320 0 8 32 0 0 5
433 613
433 750
945 750
945 722
955 722
1 1 5 0 0 8320 0 24 6 0 0 4
725 720
725 652
411 652
411 613
1 1 6 0 0 8320 0 5 25 0 0 4
181 628
181 670
781 670
781 669
0 1 7 0 0 4096 0 0 12 7 0 3
107 671
107 725
110 725
1 1 8 0 0 8320 0 2 10 0 0 7
365 613
365 654
98 654
98 761
98 761
98 758
108 758
1 1 7 0 0 20624 0 1 9 0 0 7
132 630
132 671
107 671
107 671
153 671
153 740
161 740
1 1 9 0 0 16512 0 17 3 0 0 5
348 743
337 743
337 716
388 716
388 613
1 1 10 0 0 8320 0 4 16 0 0 3
157 631
157 708
434 708
3 1 11 0 0 8320 0 34 38 0 0 3
1125 786
1169 786
1169 610
3 1 12 0 0 8320 0 29 37 0 0 3
1125 734
1137 734
1137 610
2 0 13 0 0 4224 0 29 0 0 20 2
1079 743
929 743
4 1 14 0 0 8320 0 33 29 0 0 4
1067 702
1072 702
1072 725
1079 725
2 2 15 0 0 4224 0 30 35 0 0 2
979 777
1015 777
2 3 16 0 0 16512 0 31 33 0 0 5
882 788
882 787
937 787
937 711
1022 711
0 1 17 0 0 4096 0 0 31 18 0 3
843 811
843 788
846 788
2 2 18 0 0 12416 0 32 33 0 0 4
991 722
993 722
993 702
1022 702
3 2 17 0 0 12416 0 26 34 0 0 4
829 811
863 811
863 795
1079 795
4 1 19 0 0 4224 0 35 34 0 0 2
1060 777
1079 777
3 1 13 0 0 0 0 21 30 0 0 4
917 722
929 722
929 777
943 777
2 1 20 0 0 8320 0 36 35 0 0 4
991 674
1007 674
1007 768
1015 768
0 1 3 0 0 0 0 0 36 1 0 3
950 694
950 674
955 674
0 3 4 0 0 0 0 0 35 2 0 5
945 733
945 736
980 736
980 786
1015 786
2 0 21 0 0 4224 0 21 0 0 32 2
871 731
578 731
4 1 22 0 0 8320 0 25 21 0 0 4
826 678
836 678
836 713
871 713
2 2 23 0 0 4224 0 22 27 0 0 2
634 770
726 770
2 3 24 0 0 12416 0 23 25 0 0 4
593 787
661 787
661 687
781 687
0 1 25 0 0 4096 0 0 23 30 0 3
549 807
549 787
557 787
2 2 26 0 0 8320 0 24 25 0 0 4
761 720
769 720
769 678
781 678
3 2 25 0 0 12416 0 15 26 0 0 6
529 807
557 807
557 806
728 806
728 820
783 820
4 1 27 0 0 4224 0 27 26 0 0 3
771 770
771 802
783 802
3 1 21 0 0 0 0 20 22 0 0 6
550 726
550 725
578 725
578 771
598 771
598 770
2 1 28 0 0 12416 0 28 27 0 0 4
610 695
647 695
647 761
726 761
0 1 6 0 0 0 0 0 28 4 0 3
183 670
574 670
574 695
0 3 5 0 0 0 0 0 27 3 0 3
706 652
706 779
726 779
2 0 29 0 0 12416 0 20 0 0 44 4
504 735
478 735
478 757
217 757
4 1 30 0 0 4224 0 16 20 0 0 2
479 717
504 717
2 2 31 0 0 8320 0 19 14 0 0 3
308 770
308 774
429 774
2 3 32 0 0 4224 0 18 16 0 0 4
285 799
407 799
407 726
434 726
0 1 33 0 0 4096 0 0 18 42 0 3
226 798
249 798
249 799
2 2 34 0 0 12416 0 17 16 0 0 4
384 743
400 743
400 717
434 717
3 2 33 0 0 12416 0 11 15 0 0 4
211 798
226 798
226 816
483 816
4 1 35 0 0 4224 0 14 15 0 0 3
474 774
474 798
483 798
3 1 29 0 0 0 0 9 19 0 0 4
206 749
217 749
217 770
272 770
2 1 36 0 0 8320 0 13 14 0 0 4
378 688
381 688
381 765
429 765
0 1 10 0 0 0 0 0 13 9 0 3
332 708
332 688
342 688
0 3 9 0 0 0 0 0 14 8 0 3
337 716
337 783
429 783
2 2 37 0 0 8320 0 12 11 0 0 4
146 725
147 725
147 807
166 807
0 1 8 0 0 0 0 0 11 6 0 3
98 761
98 789
166 789
2 2 38 0 0 4224 0 10 9 0 0 2
144 758
161 758
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 122
53 476 400 540
64 484 388 532
122 b) Implementamos um circuito l�gico que retorna X=1 se 
o n�mero A: (A3A2A1A0) > B: (B3B2B1B0), e retorna Y=1 
se B>A.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
